library verilog;
use verilog.vl_types.all;
entity ds_types_sv_unit is
end ds_types_sv_unit;
