library verilog;
use verilog.vl_types.all;
entity ds_mon_sv_unit is
end ds_mon_sv_unit;
