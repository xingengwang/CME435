parameter DS_BUS_WIDTH = 8;

typedef logic [DS_BUS_WIDTH-1:0] ds_data_t;

