// NOTHING MORE TO DO HERE FOR LAB 4
parameter IN_BUS_WIDTH = 8;

typedef logic [IN_BUS_WIDTH-1:0] in_data_t;

