library verilog;
use verilog.vl_types.all;
entity ds_drvr_sv_unit is
end ds_drvr_sv_unit;
