library verilog;
use verilog.vl_types.all;
entity us_drvr_sv_unit is
end us_drvr_sv_unit;
