// NOTHING MORE TO DO HERE FOR THE LAB
parameter IN_BUS_WIDTH = 8;

typedef logic [IN_BUS_WIDTH-1:0] in_data_t;

