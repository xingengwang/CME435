library verilog;
use verilog.vl_types.all;
entity env_m is
end env_m;
