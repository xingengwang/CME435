module Program_Memory_ROM (
	input logic clock,
	input logic [7:0] address,
	output logic [7:0] q
	);

logic [7:0] ROM_Data [0:255] = '{
	8'H50,	// 00		LOAD M, #4'H00
	8'HE1,	// 01		JMP	LOOPIPINS
	8'H00,	// 02			
	8'H00,	// 03			
	8'H00,	// 04			
	8'H00,	// 05			
	8'H00,	// 06			
	8'H00,	// 07			
	8'H00,	// 08			
	8'H00,	// 09			
	8'H00,	// 0A			
	8'H00,	// 0B			
	8'H00,	// 0C			
	8'H00,	// 0D			
	8'H00,	// 0E			
	8'H00,	// 0F			
	8'HB6,	// 10	LOOPIPINS:	LOOPIPINS:	MOV I, IPINS
	8'HBF,	// 11		MOV dm, IPINS
	8'HA7,	// 12		MOV OREG, dm
	8'HE1,	// 13		JMP	LOOPIPINS
	8'H00,	// 14			
	8'H00,	// 15			
	8'H00,	// 16			
	8'H00,	// 17			
	8'H00,	// 18			
	8'H00,	// 19			
	8'H00,	// 1A			
	8'H00,	// 1B			
	8'H00,	// 1C			
	8'H00,	// 1D			
	8'H00,	// 1E			
	8'H00,	// 1F			
	8'H00,	// 20			
	8'H00,	// 21			
	8'H00,	// 22			
	8'H00,	// 23			
	8'H00,	// 24			
	8'H00,	// 25			
	8'H00,	// 26			
	8'H00,	// 27			
	8'H00,	// 28			
	8'H00,	// 29			
	8'H00,	// 2A			
	8'H00,	// 2B			
	8'H00,	// 2C			
	8'H00,	// 2D			
	8'H00,	// 2E			
	8'H00,	// 2F			
	8'H00,	// 30			
	8'H00,	// 31			
	8'H00,	// 32			
	8'H00,	// 33			
	8'H00,	// 34			
	8'H00,	// 35			
	8'H00,	// 36			
	8'H00,	// 37			
	8'H00,	// 38			
	8'H00,	// 39			
	8'H00,	// 3A			
	8'H00,	// 3B			
	8'H00,	// 3C			
	8'H00,	// 3D			
	8'H00,	// 3E			
	8'H00,	// 3F			
	8'H00,	// 40			
	8'H00,	// 41			
	8'H00,	// 42			
	8'H00,	// 43			
	8'H00,	// 44			
	8'H00,	// 45			
	8'H00,	// 46			
	8'H00,	// 47			
	8'H00,	// 48			
	8'H00,	// 49			
	8'H00,	// 4A			
	8'H00,	// 4B			
	8'H00,	// 4C			
	8'H00,	// 4D			
	8'H00,	// 4E			
	8'H00,	// 4F			
	8'H00,	// 50			
	8'H00,	// 51			
	8'H00,	// 52			
	8'H00,	// 53			
	8'H00,	// 54			
	8'H00,	// 55			
	8'H00,	// 56			
	8'H00,	// 57			
	8'H00,	// 58			
	8'H00,	// 59			
	8'H00,	// 5A			
	8'H00,	// 5B			
	8'H00,	// 5C			
	8'H00,	// 5D			
	8'H00,	// 5E			
	8'H00,	// 5F			
	8'H00,	// 60			
	8'H00,	// 61			
	8'H00,	// 62			
	8'H00,	// 63			
	8'H00,	// 64			
	8'H00,	// 65			
	8'H00,	// 66			
	8'H00,	// 67			
	8'H00,	// 68			
	8'H00,	// 69			
	8'H00,	// 6A			
	8'H00,	// 6B			
	8'H00,	// 6C			
	8'H00,	// 6D			
	8'H00,	// 6E			
	8'H00,	// 6F			
	8'H00,	// 70			
	8'H00,	// 71			
	8'H00,	// 72			
	8'H00,	// 73			
	8'H00,	// 74			
	8'H00,	// 75			
	8'H00,	// 76			
	8'H00,	// 77			
	8'H00,	// 78			
	8'H00,	// 79			
	8'H00,	// 7A			
	8'H00,	// 7B			
	8'H00,	// 7C			
	8'H00,	// 7D			
	8'H00,	// 7E			
	8'H00,	// 7F			
	8'H00,	// 80			
	8'H00,	// 81			
	8'H00,	// 82			
	8'H00,	// 83			
	8'H00,	// 84			
	8'H00,	// 85			
	8'H00,	// 86			
	8'H00,	// 87			
	8'H00,	// 88			
	8'H00,	// 89			
	8'H00,	// 8A			
	8'H00,	// 8B			
	8'H00,	// 8C			
	8'H00,	// 8D			
	8'H00,	// 8E			
	8'H00,	// 8F			
	8'H00,	// 90			
	8'H00,	// 91			
	8'H00,	// 92			
	8'H00,	// 93			
	8'H00,	// 94			
	8'H00,	// 95			
	8'H00,	// 96			
	8'H00,	// 97			
	8'H00,	// 98			
	8'H00,	// 99			
	8'H00,	// 9A			
	8'H00,	// 9B			
	8'H00,	// 9C			
	8'H00,	// 9D			
	8'H00,	// 9E			
	8'H00,	// 9F			
	8'H00,	// A0			
	8'H00,	// A1			
	8'H00,	// A2			
	8'H00,	// A3			
	8'H00,	// A4			
	8'H00,	// A5			
	8'H00,	// A6			
	8'H00,	// A7			
	8'H00,	// A8			
	8'H00,	// A9			
	8'H00,	// AA			
	8'H00,	// AB			
	8'H00,	// AC			
	8'H00,	// AD			
	8'H00,	// AE			
	8'H00,	// AF			
	8'H00,	// B0			
	8'H00,	// B1			
	8'H00,	// B2			
	8'H00,	// B3			
	8'H00,	// B4			
	8'H00,	// B5			
	8'H00,	// B6			
	8'H00,	// B7			
	8'H00,	// B8			
	8'H00,	// B9			
	8'H00,	// BA			
	8'H00,	// BB			
	8'H00,	// BC			
	8'H00,	// BD			
	8'H00,	// BE			
	8'H00,	// BF			
	8'H00,	// C0			
	8'H00,	// C1			
	8'H00,	// C2			
	8'H00,	// C3			
	8'H00,	// C4			
	8'H00,	// C5			
	8'H00,	// C6			
	8'H00,	// C7			
	8'H00,	// C8			
	8'H00,	// C9			
	8'H00,	// CA			
	8'H00,	// CB			
	8'H00,	// CC			
	8'H00,	// CD			
	8'H00,	// CE			
	8'H00,	// CF			
	8'H00,	// D0			
	8'H00,	// D1			
	8'H00,	// D2			
	8'H00,	// D3			
	8'H00,	// D4			
	8'H00,	// D5			
	8'H00,	// D6			
	8'H00,	// D7			
	8'H00,	// D8			
	8'H00,	// D9			
	8'H00,	// DA			
	8'H00,	// DB			
	8'H00,	// DC			
	8'H00,	// DD			
	8'H00,	// DE			
	8'H00,	// DF			
	8'H00,	// E0			
	8'H00,	// E1			
	8'H00,	// E2			
	8'H00,	// E3			
	8'H00,	// E4			
	8'H00,	// E5			
	8'H00,	// E6			
	8'H00,	// E7			
	8'H00,	// E8			
	8'H00,	// E9			
	8'H00,	// EA			
	8'H00,	// EB			
	8'H00,	// EC			
	8'H00,	// ED			
	8'H00,	// EE			
	8'H00,	// EF			
	8'H00,	// F0			
	8'H00,	// F1			
	8'H00,	// F2			
	8'H00,	// F3			
	8'H00,	// F4			
	8'H00,	// F5			
	8'H00,	// F6			
	8'H00,	// F7			
	8'H00,	// F8			
	8'H00,	// F9			
	8'H00,	// FA			
	8'H00,	// FB			
	8'H00,	// FC			
	8'H00,	// FD			
	8'H00,	// FE			
	8'H00 	// FF			
	};

	always @ (posedge clock)
		q <= ROM_Data[address];

endmodule
