// Global environment and test program settings

`timescale	1ns/1ns					// time units/time precision
`define		CLOCK_CYCLE 1000	// 1000 * time units = 1MHz
