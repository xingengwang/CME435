library verilog;
use verilog.vl_types.all;
entity sanity_test_p is
end sanity_test_p;
