library verilog;
use verilog.vl_types.all;
entity sanity_test is
end sanity_test;
