// TO DO: Define any constants and types that will assist
//        with the implementation of the output interface
//		    or monitor.
