// TO DO: Define any constants and types that will assist
//        with the implementation of the input interface
//		    or driver.


