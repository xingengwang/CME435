parameter OUT_LEN_BUS_WIDTH  = 5;
parameter OUT_DATA_BUS_WIDTH = 8;

typedef logic [OUT_LEN_BUS_WIDTH-1:0]  out_len_t;
typedef logic [OUT_DATA_BUS_WIDTH-1:0] out_data_t;

