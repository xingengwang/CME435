// Define any global definitions needed in the env.sv and test.sv

`timescale 1ns/1ns
`define CLOCK_CYCLE 1000
