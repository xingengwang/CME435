library verilog;
use verilog.vl_types.all;
entity us_types_sv_unit is
end us_types_sv_unit;
