library verilog;
use verilog.vl_types.all;
entity sanity_test_sv_unit is
end sanity_test_sv_unit;
