library verilog;
use verilog.vl_types.all;
entity env_sv_unit is
end env_sv_unit;
