library verilog;
use verilog.vl_types.all;
entity us_mon_sv_unit is
end us_mon_sv_unit;
