// TO DO: Define any constants and types that will assist
//        with the implementation of the input intrerface
//		  or driver.


